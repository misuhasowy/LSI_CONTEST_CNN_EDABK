
defparam AESL_inst_encode.conv1_out_U.DEPTH = 2'd2;
defparam AESL_inst_encode.pool1_out_U.DEPTH = 2'd2;
defparam AESL_inst_encode.conv2_out_U.DEPTH = 2'd2;
defparam AESL_inst_encode.pool2_out_U.DEPTH = 2'd2;
defparam AESL_inst_encode.conv3_out_U.DEPTH = 2'd2;
