
defparam AESL_inst_decode.conv4_out_U.DEPTH = 2'd2;
defparam AESL_inst_decode.upsamp4_out_U.DEPTH = 2'd2;
defparam AESL_inst_decode.conv5_out_U.DEPTH = 2'd2;
defparam AESL_inst_decode.upsamp5_out_U.DEPTH = 2'd2;
defparam AESL_inst_decode.conv6_out_U.DEPTH = 2'd2;
defparam AESL_inst_decode.upsamp6_out_U.DEPTH = 2'd2;
